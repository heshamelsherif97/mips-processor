module cpu (clk, reset);

input clk, reset;



endmodule


