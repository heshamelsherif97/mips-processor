module mips_project(input i1, output out);
assign out=i1&i1;
endmodule